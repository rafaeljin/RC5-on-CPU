LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; --use CONV_INTEGER

ENTITY IM IS
PORT(
	pc: in std_logic_vector(31 downto 0);
	inst: out STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END IM;

ARCHITECTURE Behavioral OF IM IS
	TYPE myarray IS ARRAY (0 TO 700) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	signal inst_memory: myarray:=(
"00101000","00011011","00000000","00000110",
"00000111","01111011","11111111","11111111",
"00000011","01001010","10101000","00010010",
"00000011","01011010","11010000","00010000",
"00101000","00010101","00000000","00000001",
"00000111","01011010","00000000","00000001",
"00101000","00000000","11111111","11111001",
"00101111","00001010","00000000","00000001",
"00110000","00000000","00000000","00110100",
"00101111","00001011","00000000","00000001",
"00110000","00000000","00000000","00111101",
"00101111","00001100","00000000","00000001",
"00110000","00000000","00000000","01011010",
"00101111","00001101","00000000","00000001",
"00110000","00000000","00000000","01100111",
"00101111","00001110","00000000","00000001",
"00110000","00000000","00000000","01111011",
"00110000","00000000","00000000","10001010",
"00010000","00010000","00000000","00010000",
"00010000","00001010","10000000","00000000",
"00010000","00001011","10110111","11100001",
"00010000","00001100","10011110","00110111",
"00000110","00010000","11111111","11111111",
"00000001","01001010","01010000","00010000",
"00000001","01101011","01011000","00010000",
"00000001","10001100","01100000","00010000",
"00101100","00010000","11111111","11111011",
"00000101","01101011","01010001","01100011",
"00000101","10001100","01111001","10111001",
"00000100","00001101","00000000","00000000",
"00000101","10101110","00000000","01101000",
"00000101","11001111","00000000","00010000",
"00000000","00001011","00110000","00010000",
"00000000","00001101","00101000","00010000",
"00000101","10100111","00000000","01100100",
"00100000","10100110","00000000","00000000",
"00000100","10100101","00000000","00000100",
"00000000","11001100","00110000","00010000",
"00100000","10100110","00000000","00000000",
"00101100","10100111","11111111","11111100",
"00000101","10100101","00000000","00000000",
"00000101","11001000","00000000","00000000",
"00000000","00000000","00110000","00010000",
"00000000","00000000","01001000","00010000",
"00000100","00000111","00000000","01001110",
"00000001","00100110","00110000","00010000",
"00011100","10100010","00000000","00000000",
"00000000","01000110","00110000","00010000",
"00010000","00011011","00000000","00000011",
"00000000","00000110","11010000","00010011",
"00000000","00001010","11000000","00010011",
"00110000","00000000","00000000","00000000",
"00000111","01000110","00000000","00000000",
"00100000","10100110","00000000","00000000",
"00000001","00100110","01001000","00010000",
"00001101","00111011","00000000","00011111",
"00011101","00000010","00000000","00000000",
"00000001","00100010","01001000","00010000",
"00000000","00001001","11010000","00010011",
"00000000","00001011","11000000","00010011",
"00110000","00000000","00000000","00000000",
"00000111","01001001","00000000","00000000",
"00100001","00001001","00000000","00000000",
"00000100","10100101","00000000","00000100",
"00101100","10101110","00000000","00000001",
"00000111","10100101","00000000","00000000",
"00000101","00001000","00000000","00000100",
"00101101","00001111","00000000","00000001",
"00000101","11001000","00000000","00000000",
"00000100","11100111","11111111","11111111",
"00101100","00000111","11111111","11100110",
"00011101","11100010","00000000","00000000",
"00011101","11100011","00000000","00000100",
"00101100","00011111","00000000","00100110",
"00000101","10100101","00000000","00000000",
"00011100","10100110","00000000","00000000",
"00000000","01000110","00010000","00010000",
"00000100","10100101","00000000","00000100",
"00011100","10100110","00000000","00000000",
"00000000","01100110","00011000","00010000",
"00000100","00001001","00000000","00001100",
"00000000","00000010","10110000","00010100",
"00000000","00000011","10111000","00010100",
"00000000","01000011","00010000","00010011",
"00000010","11010111","10110000","00010011",
"00000000","01010110","00010000","00010010",
"00001100","01111011","00000000","00011111",
"00000000","00000010","11010000","00010011",
"00000000","00001100","11000000","00010011",
"00110000","00000000","00000000","00000000",
"00000111","01000010","00000000","00000000",
"00000100","10100101","00000000","00000100",
"00011100","10100110","00000000","00000000",
"00000000","01000110","00010000","00010000",
"00011101","11111111","00000000","00001000",
"00000000","00000010","10110000","00010100",
"00000000","01000011","00011000","00010011",
"00000010","11010111","10111000","00010011",
"00000000","01110111","00011000","00010010",
"00001100","01011011","00000000","00011111",
"00000000","00000011","11010000","00010011",
"00000000","00001101","11000000","00010011",
"00110000","00000000","00000000","00000000",
"00000111","01000011","00000000","00000000",
"00000100","10100101","00000000","00000100",
"00011100","10100110","00000000","00000000",
"00000000","01100110","00011000","00010000",
"00000101","00101001","11111111","11111111",
"00101101","00100000","11111111","11100100",
"00100001","11100011","00000000","00000100",
"00100001","11100010","00000000","00000000",
"11111111","11111111","11111111","11111111",
"00000101","11000101","00000000","00000000",
"00000100","00001001","00000000","00001100",
"00001000","10100101","00000000","00000100",
"00011100","10100110","00000000","00000000",
"00000000","01100110","00011000","00010001",
"00000000","00000010","10110000","00010100",
"00000110","11010110","00000000","00000001",
"00001110","11011011","00000000","00011111",
"00000000","00000011","11010000","00010011",
"00000000","00001110","11000000","00010011",
"00110000","00000000","00000000","00000000",
"00000111","01000011","00000000","00000000",
"00000000","00000011","10111000","00010100",
"00000000","00000010","10110000","00010100",
"00000000","01000011","00011000","00010011",
"00000010","11010111","10111000","00010011",
"00000000","01110111","00011000","00010010",
"00001000","10100101","00000000","00000100",
"00011100","10100110","00000000","00000000",
"00000000","01000110","00010000","00010001",
"00000000","00000011","10111000","00010100",
"00000110","11110111","00000000","00000001",
"00001110","11111011","00000000","00011111",
"00000000","00000010","11010000","00010011",
"00000000","00001111","11000000","00010011",
"00110000","00000000","00000000","00000000",
"00000111","01000010","00000000","00000000",
"00000000","00000010","10110000","00010100",
"00000000","00000011","10111000","00010100",
"00000000","01000011","00010000","00010011",
"00000010","11010111","10110000","00010011",
"00000000","01010110","00010000","00010010",
"00000101","00101001","11111111","11111111",
"00101100","00001001","11111111","11100000",
"00011101","10100110","00000000","00000100",
"00000000","01100110","00011000","00010001",
"00011101","10100110","00000000","00000000",
"00000000","01000110","00010000","00010001",
"00100001","11100011","00000000","00000100",
"00100001","11100010","00000000","00000000",
"11111111","11111111","11111111","11111111",
"00000000","00000000","00000000","00000000",
-- write to reg31 
"00011100","00011111","00000000","10000000",
"00110000","00000000","00000000","00010010",
		others=>(others=>'0'));
		
	attribute ram_style: string;
	attribute ram_style of inst_memory : signal is "block";
BEGIN
	-- pc(8 downto 0)?
	inst <= 	inst_memory(CONV_INTEGER(pc)) & 
				inst_memory(CONV_INTEGER(pc)+1) & 
				inst_memory(CONV_INTEGER(pc)+2) & 
				inst_memory(CONV_INTEGER(pc)+3);
END Behavioral;